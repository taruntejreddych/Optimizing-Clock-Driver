magic
tech scmos
timestamp 1574435001
<< nwell >>
rect 91 59 212 226
rect -25 3 16 33
rect 26 3 76 45
rect 90 4 212 59
rect 263 5 409 1658
rect 91 3 212 4
<< ntransistor >>
rect -6 -15 -3 -11
rect 43 -29 46 -17
rect 140 -109 143 -21
<< ptransistor >>
rect -6 10 -3 19
rect 43 9 46 35
rect 140 11 143 215
<< ndiffusion >>
rect -16 -15 -13 -11
rect -9 -15 -6 -11
rect -3 -15 0 -11
rect 4 -15 8 -11
rect 34 -21 43 -17
rect 34 -25 36 -21
rect 40 -25 43 -21
rect 34 -29 43 -25
rect 46 -21 65 -17
rect 46 -25 53 -21
rect 57 -25 65 -21
rect 46 -29 65 -25
rect 94 -48 140 -21
rect 94 -52 100 -48
rect 104 -52 140 -48
rect 94 -109 140 -52
rect 143 -47 197 -21
rect 143 -51 156 -47
rect 160 -51 197 -47
rect 143 -109 197 -51
rect 282 -78 401 -63
rect 282 -82 380 -78
rect 384 -82 401 -78
rect 282 -164 401 -82
rect 282 -168 285 -164
rect 289 -168 401 -164
rect 282 -751 401 -168
<< pdiffusion >>
rect 274 252 398 1639
rect 274 248 282 252
rect 286 248 398 252
rect 101 90 140 215
rect 101 85 106 90
rect 110 85 140 90
rect 33 24 43 35
rect 33 20 37 24
rect 41 20 43 24
rect -16 17 -6 19
rect -16 13 -14 17
rect -10 13 -6 17
rect -16 10 -6 13
rect -3 17 6 19
rect -3 13 0 17
rect 4 13 6 17
rect -3 10 6 13
rect 33 9 43 20
rect 46 23 64 35
rect 46 19 53 23
rect 57 19 64 23
rect 46 9 64 19
rect 101 11 140 85
rect 143 26 188 215
rect 143 22 156 26
rect 160 22 188 26
rect 143 11 188 22
rect 274 36 398 248
rect 274 32 380 36
rect 384 32 398 36
rect 274 20 398 32
<< ndcontact >>
rect -13 -15 -9 -11
rect 0 -15 4 -11
rect 36 -25 40 -21
rect 53 -25 57 -21
rect -13 -43 -9 -39
rect 100 -52 104 -48
rect -13 -66 -9 -61
rect 36 -67 40 -63
rect -13 -100 -9 -95
rect 36 -99 40 -95
rect 156 -51 160 -47
rect 380 -82 384 -78
rect 100 -124 104 -120
rect -13 -133 -9 -128
rect 36 -133 40 -129
rect 100 -146 104 -142
rect -13 -168 -9 -164
rect 36 -168 40 -164
rect 100 -168 104 -164
rect 285 -168 289 -164
<< pdcontact >>
rect -14 248 -10 252
rect 37 248 41 252
rect 106 248 110 252
rect 152 248 156 252
rect 219 248 223 252
rect 282 248 286 252
rect 37 207 41 211
rect -14 200 -10 204
rect -14 167 -10 171
rect 37 168 41 172
rect -14 119 -10 123
rect 37 122 41 126
rect 106 85 110 90
rect -14 66 -10 70
rect 37 68 41 72
rect 37 20 41 24
rect -14 13 -10 17
rect 0 13 4 17
rect 53 19 57 23
rect 156 22 160 26
rect 380 32 384 36
<< polysilicon >>
rect 140 215 143 231
rect -6 19 -3 39
rect 43 35 46 49
rect -6 -11 -3 10
rect -6 -19 -3 -15
rect 43 -17 46 9
rect 140 -21 143 11
rect 43 -40 46 -29
rect 140 -123 143 -109
<< polycontact >>
rect -12 -5 -6 0
rect 37 -6 43 -1
rect 134 -7 140 -1
rect 373 -7 380 -1
<< metal1 >>
rect -10 248 37 252
rect 41 248 106 252
rect 110 248 152 252
rect 156 248 219 252
rect 223 248 282 252
rect -14 204 -10 248
rect -14 171 -10 200
rect -14 123 -10 167
rect -14 70 -10 119
rect -14 17 -10 66
rect 37 211 41 248
rect 37 172 41 207
rect 37 126 41 168
rect 37 72 41 122
rect 106 90 110 248
rect 37 24 41 68
rect -43 -5 -12 0
rect 0 -1 4 13
rect 53 -1 57 19
rect 156 -1 160 22
rect 0 -6 37 -1
rect 0 -11 4 -6
rect 53 -7 134 -1
rect 156 -7 373 -1
rect -13 -39 -9 -15
rect 53 -21 57 -7
rect -13 -61 -9 -43
rect -13 -95 -9 -66
rect -13 -128 -9 -100
rect -13 -164 -9 -133
rect 36 -63 40 -25
rect 156 -47 160 -7
rect 36 -95 40 -67
rect 36 -129 40 -99
rect 36 -164 40 -133
rect 380 -15 384 32
rect 380 -22 465 -15
rect 100 -120 104 -52
rect 380 -78 384 -22
rect 100 -142 104 -124
rect 100 -164 104 -146
rect -9 -168 36 -164
rect 40 -168 100 -164
rect 104 -168 285 -164
<< labels >>
rlabel metal1 13 -166 13 -166 1 gnd
rlabel metal1 1 250 1 250 1 vdd
rlabel metal1 -26 -2 -26 -2 1 vin
rlabel metal1 449 -18 449 -18 1 vout
<< end >>
